
module toy_mem_adapter #(

) (
    input       clk         ,
    input       rst_n       ,

    

);

endmodule